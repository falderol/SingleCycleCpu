LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE work.reg_type.all;

ENTITY test_bench_Dec_5x32 IS
END test_bench_Dec_5x32;

ARCHITECTURE test OF test_bench_Dec_5x32 IS
    SIGNAL testInput: reg_address;
    SIGNAL testEnable: STD_LOGIC; 
    SIGNAL testOutput: STD_LOGIC_VECTOR(31 DOWNTO 0);

BEGIN
    test5x32: ENTITY work.DEC_5x32(logic) PORT MAP (testInput, testEnable, testOutput);
    PROCESS
    TYPE pattern_type IS RECORD
        Input_5x32: reg_address;
        Enable_5x32: STD_LOGIC;
        Output_5x32: STD_LOGIC_VECTOR(31 DOWNTO 0);
    END RECORD;

    TYPE pattern_array IS ARRAY (NATURAL RANGE <>) OF pattern_type;
        CONSTANT patterns: pattern_array :=
            ( ("00000", '1', "00000000000000000000000000000001"),
              ("00001", '1', "00000000000000000000000000000010"),
              ("00010", '1', "00000000000000000000000000000100"),
              ("00011", '1', "00000000000000000000000000001000"),
              ("00100", '1', "00000000000000000000000000010000"),
              ("00101", '1', "00000000000000000000000000100000"),
              ("00110", '1', "00000000000000000000000001000000"),
              ("00111", '1', "00000000000000000000000010000000"),
              ("01000", '1', "00000000000000000000000100000000"),
              ("01001", '1', "00000000000000000000001000000000"),
              ("01010", '1', "00000000000000000000010000000000"),
              ("01011", '1', "00000000000000000000100000000000"),
              ("01100", '1', "00000000000000000001000000000000"),
              ("01101", '1', "00000000000000000010000000000000"),
              ("01110", '1', "00000000000000000100000000000000"),
              ("01111", '1', "00000000000000001000000000000000"),
              ("10000", '1', "00000000000000010000000000000000"),
              ("10001", '1', "00000000000000100000000000000000"),
              ("10010", '1', "00000000000001000000000000000000"),
              ("10011", '1', "00000000000010000000000000000000"),
              ("10100", '1', "00000000000100000000000000000000"),
              ("10101", '1', "00000000001000000000000000000000"),
              ("10110", '1', "00000000010000000000000000000000"),
              ("10111", '1', "00000000100000000000000000000000"),
              ("11000", '1', "00000001000000000000000000000000"),
              ("11001", '1', "00000010000000000000000000000000"),
              ("11010", '1', "00000100000000000000000000000000"),
              ("11011", '1', "00001000000000000000000000000000"),
              ("11100", '1', "00010000000000000000000000000000"),
              ("11101", '1', "00100000000000000000000000000000"),
              ("11110", '1', "01000000000000000000000000000000"),
              ("11111", '1', "10000000000000000000000000000000"),
              ("11111", '0', "00000000000000000000000000000000")
            );
    BEGIN
        FOR i In patterns'range LOOP
            testInput <= patterns(i).Input_5x32;
            testEnable <= patterns(i).Enable_5x32;
        wait for 1 ms;
 
        assert testOutput = patterns(i).Output_5x32
            report "bad output" severity error;
        END LOOP;

        assert false
            report "end of test" severity note;
        wait;
    END PROCESS;
END test;


