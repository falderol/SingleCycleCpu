LIBRARY ieee;
USE ieee.std_logic_1164.all;

PACKAGE op_type IS 
    SUBTYPE op IS STD_LOGIC_VECTOR(3 DOWNTO 0);
END op_type;


