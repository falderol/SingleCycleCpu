LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE work.word_type.all;

ENTITY test_bench_32x32x1_vector IS
END test_bench_32x32x1_vector;

ARCHITECTURE test OF test_bench_32x32x1_vector IS
    SIGNAL testI: word_array;
    SIGNAL testS: STD_LOGIC_VECTOR(4 DOWNTO 0);
    SIGNAL testOUT: word;

BEGIN
    test32: ENTITY work.MUX_32x32x1_vector(logic) PORT MAP ( testI, testS, testOUT );
    PROCESS
        TYPE pattern_type IS RECORD
            I: word_array;
            S: STD_LOGIC_VECTOR(4 DOWNTO 0);
            o: word;
        END RECORD;

        TYPE pattern_array IS ARRAY (NATURAL RANGE <>) OF pattern_type;
        CONSTANT patterns: pattern_array :=
-- All 1's I00, All 0's I31
            ( ( ("00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000001"
               ),
                 "00000",
                 "00000000000000000000000000000001"
              ),
              ( ("00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000001",
                 "00000000000000000000000000000000"
               ),
                 "00001",
                 "00000000000000000000000000000001"
              ),

              ( ("00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000001",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000"
               ),
                 "00010",
                 "00000000000000000000000000000001"
              ),


              ( ("00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000001",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000"
               ),
                 "00100",
                 "00000000000000000000000000000001"
              ),

              ( ("00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000001",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000"
               ),
                 "01000",
                 "00000000000000000000000000000001"
              ),

              ( ("00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000001",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000"
               ),
                 "10000",
                 "00000000000000000000000000000001"
              ),

              ( ("00000000000000000000000000000001",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000",
                 "00000000000000000000000000000000"
              ),
                 "11111",
                 "00000000000000000000000000000001"
              ) 
            );
    BEGIN
        FOR i IN patterns'range LOOP
            testI <= patterns(i).I;
            testS <= patterns(i).S;

            wait for 1 ms;

            assert testOUT = patterns(i).o
                report "bad output" severity error;
        END LOOP;

        assert false
            report "end of test" severity note;
        wait;
    END PROCESS;
END test;
